
entity myOr16 is 
	port(a, b : in bit; c : out bit); 

end myOr16;