
entity myNor is 
	port(a, b : in bit; c : out bit); 

end myNor;