
entity myDMux16 is 
	port(a, b : in bit; c : out bit); 

end myDMux16;