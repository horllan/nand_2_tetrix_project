
entity myMux16 is 
	port(a, b : in bit; c : out bit); 

end myMux16;